* D:\kicad works\ajay\doorbell\door.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/28/18 11:49:36

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_P1-Pad1_ Net-_P1-Pad2_ BC547		
Q2  Net-_P2-Pad2_ Net-_Q2-Pad2_ Net-_P1-Pad2_ BC548		
P1  Net-_P1-Pad1_ Net-_P1-Pad2_ CONN_01X02		
P2  Net-_P1-Pad1_ Net-_P2-Pad2_ CONN_01X02		
R1  Net-_Q2-Pad2_ Net-_Q1-Pad1_ R		

.end
